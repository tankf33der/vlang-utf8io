module utf8io

fn test_peek() {
	u := utf8io.Utf8io{}
	unsafe { u.free() }
}
