module utf8io

fn test_to_arrays_ascii() {
	println(utf8io.to_arrays('mike'))
	assert true
}

