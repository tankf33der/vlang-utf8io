module utf8io

pub struct Utf8io{
pub mut:
	f	File
}

pub open(path string)! {


}

