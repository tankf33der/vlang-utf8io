module utf8io

fn test_peek() {

}
